** sch_path: /home/yogesh/invcprpd.sch
**.subckt invcprpd
XX1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VIN IN GND pulse(0 1.8 1n 0.3n 0.3n 5n 10n)
VSS1 VSS GND 0
VDD VDD GND 1.8
Xx0 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.58 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.lib /home/yogesh/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.save all

.control
  * 1. Run time simulation
  tran 0.1n 30n

  * 2. Measure 50% delay points (Input to Output)
  meas tran tpHL trig v(IN) val=0.9 rise=2 targ v(OUT) val=0.9 fall=2
  meas tran tpLH trig v(IN) val=0.9 fall=2 targ v(OUT) val=0.9 rise=2

   let p_inst = v(vdd) * -i(vdd)

  * 3. Calculate and display average delay
  let tp_avg = (tpHL + tpLH) / 2
  print tpHL tpLH tp_avg
  plot (p_inst)
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
